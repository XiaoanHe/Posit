module test_fpmultiplier;

timeunit 1ns; timeprecision 10ps;

logic signed [31:0] product;
logic ready;
logic signed [31:0] a;
logic clock;
logic nreset;



fpmultiplier Fp ( product, ready, a, clock, nreset );

always
  begin
         clock = 0;
    #250 clock = 1;
    #500 clock = 0;
    #250 clock = 0;
  end

// initial
//     begin
// 	nreset = 0;
//       #1000
// 	nreset = 0;
//       #1000
// 	nreset = 1;
//       #5000
// 	$finish;
//     end

  initial
    begin
	a = '0;

      // 0.7 * 0.1 gets 0.0699999928474
      // 00111101100011110101110000101000
      // #2000
	// a = 32'b0_01111110_01100110011001100110011;
      // #1500
      // a = 32'b0_01111011_10011001100110011001101;

      // // 0.2*0.1 gets 0.0199999995529651641845703125
      // // 00111100101000111101011100001010
      // #2000
	// a = 32'b0_01111100_10011001100110011001101;
      // #1500
      // a = 32'b0_01111011_10011001100110011001101;

      // // 33554435*33555435 gets 1.125933663e15
      // // 01011000100000000000000011110110
      // // 1125932924403712
      // #2000
	// a = 32'b0_100110000_0000000000000000000001;
      // #1500
      // a = 32'b0_10011000_00000000000000011111011;

      // 4.5e9*5.5e9 gets 2.475e19
      // 00111100101000111101011100001010
      #2000
	a = 32'b0_10011111_00001100001110001000110;
      #1500
      a = 32'b0_10011111_01000111110100110101100;
      
      // #2000
	// a = 32'b0_01111110_11001100110011001100110;
      // #1500
      // a = 32'b0_01111011_10011001100110011001101;

      // // 10000.7 * 10000.1 gets 100007992
      // // 01001100101111101100000000000111
      // #2000
	// a = 32'b01000110000111000100001011001101;
      // #1500
      // a = 32'b01000110000111000100000001100110;

      // // 10000.2*10000.1 gets 100002992
      // // 01001100101111101011110110010110
      // #2000
	// a = 32'b01000110000111000100000011001101;
      // #1500
      // a = 32'b01000110000111000100000001100110;

      // 20000.900390625 * 10000.1 gets 200010992
      // 0_10011010_01111101011111011001111
      // #2000
	// a = 32'b01000110100111000100000111001101;
      // #1500
      // a = 32'b01000110000111000100000001100110;
    end
	endmodule