`timescale 1ns/1ps
module floatadd_tb();
    reg clk,rst;
    reg [31:0] x,y,tmp_in1,tmp_in2,z1,z2,diff;
    wire [31:0] z;
    wire [1:0] overflow;
    
    fpadder floatadd_test(
        .clk(clk),
        .rst(rst),
        .x(x),
        .y(y),
        .z(z),
        .overflow(overflow)
    );
    always #(10) clk<=~clk;
    initial begin
        clk=0;
        rst=1'b0;
        #20 rst=1'b1;
        #1000
        x=32'b0_01111011_10011001100110011001101;   //  0.100000001490116119384765625
        y=32'b0_01111100_10011001100110011001101;   //  0.20000000298023223876953125

        // #1000
        // x=32'b0_10001111_00000000000000000001101;   //  65536.1015625
        // y=32'b0_10001111_00000000000000000011010;   //  65536.203125

        // #1000
        // x=32'b0_01111110_01100110011001100110011;   //  0.699999988079071044921875
        // y=32'b0_01111100_10011001100110011001101;   //  0.20000000298023223876953125
        // // 0.89999997615814208984375  00111111011001100110011001100110
        // #1000
        // x=32'b0_01111011_00011110101110000101000;   //  0.0699999928474
        // y=32'b0_01111001_01000111101011100001010;   //  0.0199999995529651641845703125

        #1000
        x=32'b01000110000111000100001011001101;   //  10000.7
        y=32'b01000110000111000100000011001101;   //  10000.2
        // 20000.900390625 01000110100111000100000111001101
        
        #1000
        x=32'b01001100101111101100000000000111;   //  100007992
        y=32'b01001100101111101011110110010110;   //  100002992

// //////      ASSOCIATIVITY       //////
        // x = '0;
        // y = '0;
        // #200
        // x = 32'b0_10010111_11110111100010100100000;
        // y = 32'b1_10010111_11110111100010100100000;
        // #200
        // tmp_in1 = z;
        // #100
        // x = tmp_in1;
        // y = 32'b00111111100000000000000000000000;
        // #200
        // z1 = z;
        // x = '0;
        // y = '0;
        // #1000
        // x = 32'b01001011111110111100010100100000;
        // y = 32'b00111111100000000000000000000000;
        // #200
        // tmp_in2 = z;
        // #200
        // y = 32'b11001011111110111100010100100000;
        // x = tmp_in2;
        // #200
        // z2 = z;
        // #200
        // diff = z1 - z2;
        

        // #1000    //验证下溢出 0000001E
        // x=32'h00800010;  //  1.1754965929e-38
        // y=32'h80800001;  //  1.17549449095e-38

        // #1000 //denormalized + overflow=2'b11 3f8003ff
        // x=32'h000003FF;  //1.433528329e-42
        // y=32'h3F8003FF;  //1.0001219511
        
        // #1000
        // x=32'h7F800003;
        // y=32'h7F800004;//验证NaN overflow=2'b11 FFFFFFFF
        //  #1000
        // x=32'h00000000;//
        // y=32'h9FFFFFF0;//-1.0842011385097E-19   9FFFFFF0
        // //验证判断0阶段功能
        // #1000
        // x=32'h00000003;
        // y=32'h00000005;//非规格数字+非规格 数字 00000008
        // #1000
        // x=32'h1FFFFFFF;//1.084202107862E-19
        // y=32'h9FFFFFF0;//-1.0842011385097E-19
        // //ans=0.0000009693523   15F00000
        // #1000
        // x=32'h00000003;
        // y=32'h00800002;//非规格数字+正常数字 overflow=2'b11 
        // #1000
        // x=32'h1EE2281F;//2.3945274455386E-20
        // y=32'h1FFFFFF0;//1.0842011385097E-19
        // //ans=1.32365388306356E-19 
        // #1000
        // x=32'h00000003;
        // y=32'h7F800004;//非规格数字+正常数字 overflow=2'b11 
        // #1000
        // x=32'h1EE2281F;//2.3945274455386E-20
        // y=32'h1FFFFFF0;//1.0842011385097E-19
        // //ans=1.32365388306356E-19 
        // #1000
        // x=32'h7F800000;
        // y=32'h00000003;//验证无穷大，结果为无穷大 overflow=2'b11 
        // #1000
        // x=32'h1EE2281F;//2.3945274455386E-20
        // y=32'h1FFFFFF0;//1.0842011385097E-19
        // //ans=1.32365388306356E-19 
        // #1000
        // x=32'h7F800000;
        // y=32'h1FFFFFF0;//验证无穷大，结果为无穷大 overflow=2'b11 
    end
endmodule
