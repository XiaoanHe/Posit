`timescale 1ns/1ps
module floatadd_tb();
    reg clk,rst;
    reg [31:0] x,y;
    wire [31:0] z;
    wire [1:0] overflow;
    
    fpadder floatadd_test(
        .clk(clk),
        .rst(rst),
        .x(x),
        .y(y),
        .z(z),
        .overflow(overflow)
    );
    always #(10) clk<=~clk;
    initial begin
        clk=0;
        rst=1'b0;
        #20 rst=1'b1;
        #20 x=32'b0_11011111_00000000000000000000000;//79228162514264337593543950336
        y=32'b0_11011111_00000000000000000000000;//79228162514264337593543950336
        //ans=0.78+0.55=1.33 32'b00111111 10101010 00111101 01110001 3faa3d70
        #1000   //验证上溢出 overflow=2'b01 7FFFFFFF
        x=32'h7F7FFFFF;
        y=32'h7F7FFFFF;
        #1000
        x=32'b0_00000000_00000000000000000000000;   //  0
        y=32'b0_11111110_11111111111111111111111;   //  3.40282346639e+38

        // #1000    //验证下溢出 0000001E
        // x=32'h00800010;  //  1.1754965929e-38
        // y=32'h80800001;  //  1.17549449095e-38

        // #1000 //denormalized + overflow=2'b11 3f8003ff
        // x=32'h000003FF;  //1.433528329e-42
        // y=32'h3F8003FF;  //1.0001219511
        
        // #1000
        // x=32'h7F800003;
        // y=32'h7F800004;//验证NaN overflow=2'b11 FFFFFFFF
        //  #1000
        // x=32'h00000000;//
        // y=32'h9FFFFFF0;//-1.0842011385097E-19   9FFFFFF0
        // //验证判断0阶段功能
        // #1000
        // x=32'h00000003;
        // y=32'h00000005;//非规格数字+非规格 数字 00000008
        // #1000
        // x=32'h1FFFFFFF;//1.084202107862E-19
        // y=32'h9FFFFFF0;//-1.0842011385097E-19
        // //ans=0.0000009693523   15F00000
        // #1000
        // x=32'h00000003;
        // y=32'h00800002;//非规格数字+正常数字 overflow=2'b11 
        // #1000
        // x=32'h1EE2281F;//2.3945274455386E-20
        // y=32'h1FFFFFF0;//1.0842011385097E-19
        // //ans=1.32365388306356E-19 
        // #1000
        // x=32'h00000003;
        // y=32'h7F800004;//非规格数字+正常数字 overflow=2'b11 
        // #1000
        // x=32'h1EE2281F;//2.3945274455386E-20
        // y=32'h1FFFFFF0;//1.0842011385097E-19
        // //ans=1.32365388306356E-19 
        // #1000
        // x=32'h7F800000;
        // y=32'h00000003;//验证无穷大，结果为无穷大 overflow=2'b11 
        // #1000
        // x=32'h1EE2281F;//2.3945274455386E-20
        // y=32'h1FFFFFF0;//1.0842011385097E-19
        // //ans=1.32365388306356E-19 
        // #1000
        // x=32'h7F800000;
        // y=32'h1FFFFFF0;//验证无穷大，结果为无穷大 overflow=2'b11 
        #2000 $stop;
    end
endmodule
