/////////////////////////////////////////////////////////////////////
// Design unit: Posit Adder Testbench
//            :
// File name  : Posit_Adder_32bits_tb-4.sv
//            :
// Description: Test Posit Adder
//            :
// Limitations: None
//            : 
// System     : SystemVerilog IEEE 1800-2005
//            :
// Author     : Xiaoan(Jasper) He 
//            : xh2g20@ecs.soton.ac.uk
//
// Revision   : Version 1.0 20/02/2023
/////////////////////////////////////////////////////////////////////

timeunit 1ns; timeprecision 1ps;

module Posit_Adder_32Bit_es4_tb;
parameter N = 32, RS = $clog2(N), ES = 4;

//input logic
logic signed [N-1:0] IN1, IN2, tmp_in1, tmp_in2, OUT1,OUT2,diff;

//output logic
logic signed [N-1:0] OUT;

reg clk;
bit [N-1:0]outf [100];
integer outfile;
reg start;
reg [N-1:0] data1 [1:100];
reg [N-1:0] data2 [1:100];

initial $readmemb("IN1_k=3.txt",data1);
initial $readmemb("IN2_k=3.txt",data2);
Posit_Adder #(.N(N), .ES(ES)) PA_tb (.*);
initial 
    begin
        #10
        IN1 = '0;
        IN2 = '0;

        // //////      CORNER CASES        //////
        // #90 //  3.40282346639E+38   +   3.40282346639E+38
        // IN1 = 32'b01111111110000000000000000000000;
        // IN2 = 32'b01111111110000000000000000000000;
        
        // #50 //  1.401298464324817e-45   +   1.401298464324817e-45
        // IN1 = 32'b11111111111001010000000000000000;
        // IN2 = 32'b11111111111001010000000000000000;

        // #50 //  0.7+0.2
        // IN1 = 32'b00111000001111010111000010100100;
        // IN2 = 32'b00111011001100110011001100110011;

        // #50 //  0.07+0.02
        // IN1 = 32'b00111000001111010111000010100100;
        // IN2 = 32'b00110100100011110101110000101001;

        // #50 //  90.7+85.2 = 175.9000015258789
        // IN1 = 32'b01001100110101011001100110011010;
        // IN2 = 32'b01001100101010011001100110011010;

        // #50 //  8172.072021484375 + 7676.5201416015625 = 15848.59228515625
        //     //  +1011011110111101000100101111010
        // IN1 = 32'b01011001111111011000001001001110;
        // IN2 = 32'b01011001101111111001000010100101;

        #50 //  8172.072021484375 + 7676.5201416015625 = 15848.59228515625
            //  +1011011110111101000100101111010
        IN1 = 32'b00000000000010110011111110010000;
        IN2 = 32'b00000000000010101011111110010000;
        // #50 //  10000.7+10000.2 gets 20000.89990234375
        // IN1 = 32'b01011010011100010000101100110011;
        // IN2 = 32'b01011010011100010000001100110011;

        // #50 //  100008000 + 100003000 gets 200011000
        // IN1 = 32'b01101010011111011000000000010000;
        // IN2 = 32'b01101010011111010111101100101110;

    end

    // //     //////      MIDDLE RANGE       //////
    
        
    //     reg [15:0] i;
            
    //         initial 
    //         begin
                
    //             // Initialize Inputs
    //             IN1 = 0;
    //             IN2 = 0;
    //             clk = 0;
    //             start = 0;
            
                
    //             // Wait 100 ns for global reset to finish
    //             #100 i=0;
    //             #20 start = 1;
    //                     #6000 start = 0;
    //             #100;
                
    //             $fclose(outfile);
    //             $finish;
    //         end


    //     always #5 clk=~clk;

    //     always @(posedge clk) 
    //     begin			
    //         IN1=data1[i];	
    //         IN2=data2[i];
    //         if(i==101)
    //         begin
    //             $finish;
    //         end
    //         else i = i + 1;
    //     end

    //     initial outfile = $fopen("OUTPUT_k=3.txt", "w");

    //     always @(negedge clk) 
    //     begin
    //         outf[i] = OUT;
    //         $fwrite(outfile, "%b\n", OUT);
    //     end

        //////      PRECISION       //////
    // initial
        // begin
        // #10
        // IN1 = '0;
        // IN2 = '0;
        // #90 //  0.1 + 0.2
        // IN1 = 32'b00111001001100110011001100110011;
        // IN2 = 32'b00111011001100110011001100110011;
        
        // #50 //  65536.1+65536.2
        // IN1 = 32'b01100000000000000000000000110011;
        // IN2 = 32'b01100000000000000000000000011010;

        // IN1 = 32'b01110000000000000000000000000010;
        // IN2 = 32'b01110000000000000000000000000100;

        // IN1 = 32'b01111000000001000011011001001100;
        // IN2 = 32'b01111000000000100100011000010100;
    //     end

        //////      ASSOCIATIVITY       //////
        // initial
        // begin
        // #10
        // IN1 = '0;
        // IN2 = '0;
        // #90
        // IN1 = 32'b01101000111101111000101001000000;
        // IN2 = 32'b10010111000010000111010111000000;
        // #20
        // tmp_in1 = OUT;
        // #80
        // IN1 = tmp_in1;
        // IN2 = 32'b01000000000000000000000000000000;
        // #20
        // OUT1 = OUT;
        // #100
        // IN1 = 32'b01101000111101111000101001000000; 
        // IN2 = 32'b01000000000000000000000000000000;
        // #20
        // tmp_in2 = OUT;
        // #80
        // IN1 = 32'b10010111000010000111010111000000;
        // IN2 = tmp_in2;
        // #20
        // OUT2 = OUT;
        // #50
        // diff = OUT1 - OUT2;
        // end

        // initial
        // begin
        // #10
        // IN1 = '0;
        // IN2 = '0;
        // #90
        // IN1 = 32'b01110011000101010000001011111001;
        // IN2 = 32'b10001100111010101111110100000111;
        // #20
        // tmp_in1 = OUT;
        // #80
        // IN1 = tmp_in1;
        // IN2 = 32'b01000000000000000000000000000000;
        // #20
        // OUT1 = OUT;
        // #100
        // IN1 = 32'b01110011000101010000001011111001;
        // IN2 = 32'b01000000000000000000000000000000;
        // #20
        // tmp_in2 = OUT;
        // #80
        // IN1 = 32'b10001100111010101111110100000111;
        // IN2 = tmp_in2;
        // #20
        // OUT2 = OUT;
        // #50
        // diff = OUT1 - OUT2;
        // end

    //     #90 // test action related to infinity
    //     IN1 = 32'b10000000000000000000000000000000; // inf
    //     IN2 = 32'b10101001001010101010010001010110; // random number
    // //  OUT = 32'b10000000000000000000000000000000; // inf

    //     #50
    //     IN1 = 32'b01001001010101001010011100100010; // random number
    //     IN2 = 32'b10000000000000000000000000000000; // inf
    // //  OUT = 32'b10000000000000000000000000000000;

    //     #50 // test action related to zero
    //     IN1 = 32'b00000000000000000000000000000000; // 0
    //     IN2 = 32'b01010100101010101010010101000101; // random number
    // //  OUT = 32'b01010100101010101010010101000101;

    //     #50
    //     IN1 = 32'b01001001010101001010011100100010; // random number
    //     IN2 = 32'b00000000000000000000000000000000; // 0
    // //  OUT = 32'b01001001010101001010011100100010;

    //     #50 // +max_float_real + +max_float_real
    //     IN1 = 32'b01111111110000000000000000000000;
    //     IN2 = 32'b01111111110000000000000000000000;
    // //  OUT = 32'b01111111110000100000000000000000;

    //     #50 // (-) max_float_real + (-) max_float_real
    //     IN1 = 32'b10000000010000000000000000000000;
    //     IN2 = 32'b10000000010000000000000000000000;
    // //  OUT = 32'b10000000001111100000000000000000;

    //     #50 // +max_float_real + (-)max_float_real
    //     IN1 = 32'b01111111110000000000000000000000;
    //     IN2 = 32'b10000000010000000000000000000000;
    // //  OUT = 32'b00000000000000000000000000000000;

    //     #50 //  0.1 + 0.2
    //     IN1 = 32'b0_01_1100_1001100110011001100110011;
    //     IN2 = 32'b0_01_1101_1001100110011001100110011;

    //     #50 //  0.3 - 0.2
    //     IN1 = 32'b00111000110011001100110011001101;
    //     IN2 = 32'b11000100110011001100110011001101;

        // #50
        // IN1 = 32'b0_10_0000_0000000000000000000000000;
        // IN2 = 32'b1_10_0000_0000000000000000000000000;
        // #50ns
        // IN1 = 32'b0_10_0000_0000000000000000000000000;
        // IN2 = 32'b1_10_0000_1000000000000000000000000;
    // end



endmodule